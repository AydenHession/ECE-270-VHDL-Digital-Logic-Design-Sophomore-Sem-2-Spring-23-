begin

case (state) is
  when S0 => flag <= '0';

  when S0 => flag <= '0';

  when S0 => flag <= '1';

  when S0 => flag <= '1';

  when others => flag <= '1';

end case;
end process;

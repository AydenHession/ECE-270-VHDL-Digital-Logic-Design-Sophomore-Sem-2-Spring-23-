


    wait for clk_period*2;
        ain <= "00";
    wait for clk_period*2;
        ain <= "00";
    wait for clk_period*1;
        ain <= "00";
    wait for clk_period*1;
        ain <= "00";
    wait for clk_period*2;
        ain <= "00";
    wait for clk_period*2;
        ain <= "00";
    wait for clk_period*2;
        ain <= "00";
    wait for clk_period*2;
        ain <= "00";
    wait for clk_period*2;
        ain <= "00";
    wait for clk_period*2;
        ain <= "00";
    wait for clk_period*2;
        ain <= "00";
    wait for clk_period*2;
        ain <= "00";  
    wait for clk_period*2;
        ain <= "00";


    wait;
end process;

END;    

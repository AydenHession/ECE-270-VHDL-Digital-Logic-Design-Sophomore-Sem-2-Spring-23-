begin

    a <= "0100";
    b <= "1010";
    c <= "0";

    wait for 10 ns;
    a <= "0101";
    b <= "0111";
    c <= "0";

    wait for 10 ns;
    a <= "1010";
    b <= "0111";
    c <= "0";

    wait for 10 ns;
    a <= "1100";
    b <= "0110";
    c <= "0";

    wait for 10 ns;
    a <= "0011";
    b <= "0101";
    c <= "0";

    wait for 10 ns;
    a <= "1001";
    b <= "1000";
    c <= "0";

    wait for 10 ns;
    a <= "1110";
    b <= "0001";
    c <= "1";
